library ieee;
use ieee.std_logic_1164.all;

ENTITY BANCO_REG168 IS
    PORT(WD: IN std_logic_vector(7 DOWNTO 0);
    W, RR1, RR2: IN std_logic_vector(3 DOWNTO 0); 
    CLR, CLK, WR, EN1, EN2: IN std_logic;
    RD1, RD2: OUT std_logic_vector(7 DOWNTO 0)); 
END BANCO_REG168;


ARCHITECTURE CKT OF BANCO_REG168 IS 

COMPONENT REG8 IS
    PORT( I: IN std_logic_vector(7 DOWNTO 0);
        CLK, CLR, EN: IN std_logic;
        O: OUT std_logic_vector(7 DOWNTO 0));
END COMPONENT;

COMPONENT MUX16_8 is
	port(I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15: in std_logic_vector(7 DOWNTO 0);
		S: in std_logic_vector(3 downto 0);
        EN: IN std_logic;
		O: out std_logic_vector(7 DOWNTO 0));
END COMPONENT;

COMPONENT DEMUX16 IS
	port(I, EN: in std_logic;
		S: in std_logic_vector(3 downto 0);
		LD: out std_logic_vector(15 downto 0));
END COMPONENT;

SIGNAL LD: std_logic_vector (15 DOWNTO 0);
SIGNAL IWD, R0, R1, R2, R3, R4, R5, R6, R7, R8, R9, R10, R11, R12, R13, R14, R15: STD_LOGIC_VECTOR(7 DOWNTO 0);

BEGIN 

DEF_LD: DEMUX16 PORT MAP(WR, WR, W, LD);

DEF_REGD0: REG8 PORT MAP(WD, CLK, CLR, LD(0), R0);
DEF_REGD1: REG8 PORT MAP(WD, CLK, CLR, LD(1), R1);
DEF_REGD2: REG8 PORT MAP(WD, CLK, CLR, LD(2), R2);
DEF_REGD3: REG8 PORT MAP(WD, CLK, CLR, LD(3), R3);
DEF_REGD4: REG8 PORT MAP(WD, CLK, CLR, LD(4), R4);
DEF_REGD5: REG8 PORT MAP(WD, CLK, CLR, LD(5), R5);
DEF_REGD6: REG8 PORT MAP(WD, CLK, CLR, LD(6), R6);
DEF_REGD7: REG8 PORT MAP(WD, CLK, CLR, LD(7), R7);
DEF_REGD8: REG8 PORT MAP(WD, CLK, CLR, LD(8), R8);
DEF_REGD9: REG8 PORT MAP(WD, CLK, CLR, LD(9), R9);
DEF_REGD10: REG8 PORT MAP(WD, CLK, CLR, LD(10), R10);
DEF_REGD11: REG8 PORT MAP(WD, CLK, CLR, LD(11), R11);
DEF_REGD12: REG8 PORT MAP(WD, CLK, CLR, LD(12), R12);
DEF_REGD13: REG8 PORT MAP(WD, CLK, CLR, LD(13), R13);
DEF_REGD14: REG8 PORT MAP(WD, CLK, CLR, LD(14), R14);
DEF_REGD15: REG8 PORT MAP(WD, CLK, CLR, LD(15), R15);

DEF_RD: MUX16_8 PORT MAP(R0, R1, R2, R3, R4, R5, R6, R7, R8, R9, R10, R11, R12, R13, R14, R15, RR1, EN1, RD1);

DEF_RD2: MUX16_8 PORT MAP(R0, R1, R2, R3, R4, R5, R6, R7, R8, R9, R10, R11, R12, R13, R14, R15, RR2, EN2, RD2);

END CKT;
