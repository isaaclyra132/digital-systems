library ieee;
use ieee.std_logic_1164.all;

ENTITY T_DATA is
    PORT(IR: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    PULO, D_ADDR: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    W_ADDR, RP_ADDR, RQ_ADDR: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    IR_HLT, IR_LDR, IR_STR, IR_MOV, IR_ADD, IR_SUB, IR_AND, IR_OR, IR_NOT, IR_XOR, IR_CMP, IR_JMP, IR_JNC, IR_JC, IR_JNZ, IR_JZ: OUT STD_LOGIC);
END T_DATA;


ARCHITECTURE CKT OF T_DATA IS 

COMPONENT MUX21_4 IS
    port(A, B : in std_logic_vector(3 downto 0);
	    S : in std_logic;
        O: out std_logic_vector(3 downto 0));
END COMPONENT;

SIGNAL STR, MOV: STD_LOGIC;

BEGIN 

MUX0: MUX21_4 PORT MAP(IR(11 DOWNTO 8), IR(7 DOWNTO 4), MOV, W_ADDR);
MUX1: MUX21_4 PORT MAP(IR(7 DOWNTO 4), IR(11 DOWNTO 8), STR, RP_ADDR);

IR_HLT  <= (NOT IR(15) AND NOT IR(14) AND NOT IR(13) AND NOT IR(12));
IR_LDR  <= (NOT IR(15) AND NOT IR(14) AND NOT IR(13) AND IR(12));
STR     <= (NOT IR(15) AND NOT IR(14) AND IR(13) AND NOT IR(12));
MOV     <= (NOT IR(15) AND NOT IR(14) AND IR(13) AND IR(12));
IR_ADD  <= (NOT IR(15) AND IR(14) AND NOT IR(13) AND NOT IR(12));
IR_SUB  <= (NOT IR(15) AND IR(14) AND NOT IR(13) AND IR(12));
IR_AND  <= (NOT IR(15) AND IR(14) AND IR(13) AND NOT IR(12));
IR_OR   <= (NOT IR(15) AND IR(14) AND IR(13) AND IR(12));
IR_NOT  <= (IR(15) AND NOT IR(14) AND NOT IR(13) AND NOT IR(12));
IR_XOR  <= (IR(15) AND NOT IR(14) AND NOT IR(13) AND IR(12));
IR_CMP <= (IR(15) AND NOT IR(14) AND IR(13) AND NOT IR(12));
IR_JMP  <= (IR(15) AND NOT IR(14) AND IR(13) AND IR(12));
IR_JNC  <= (IR(15) AND IR(14) AND NOT IR(13) AND NOT IR(12));
IR_JC   <= (IR(15) AND IR(14) AND NOT IR(13) AND IR(12));
IR_JNZ  <= (IR(15) AND IR(14) AND IR(13) AND NOT IR(12));
IR_JZ   <= (IR(15) AND IR(14) AND IR(13) AND IR(12));

IR_STR <= STR;
IR_MOV <= MOV;
RQ_ADDR <= IR(3 DOWNTO 0);
PULO <= IR(7 downto 0);
D_ADDR <= IR(7 downto 0);

END CKT;