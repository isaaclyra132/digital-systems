library ieee;
use ieee.std_logic_1164.all;

ENTITY BLOCKOP IS 
    PORT(R_DATA: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
        W_ADDR, RP_ADDR, RQ_ADDR: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        ULA_SW: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
        CLK, MUX_SW, W_WR, RP_RD, RQ_RD,clr: IN STD_LOGIC;
        W_DATA, S: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
        ULA_Z, ULA_CARRY: OUT STD_LOGIC
    );
END BLOCKOP;

ARCHITECTURE CKT OF BLOCKOP IS 

COMPONENT MUX21_8 IS
	port (A, B : in STD_LOGIC_VECTOR(7 downto 0);
		S: in STD_LOGIC;
		O: out STD_LOGIC_VECTOR(7 downto 0) );
END COMPONENT;

COMPONENT BANCO_REG168 IS
    PORT(WD: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
        W, RR1, RR2: IN STD_LOGIC_VECTOR(3 DOWNTO 0); 
        CLR, CLK, WR, EN1, EN2: IN STD_LOGIC;
        RD1, RD2: OUT STD_LOGIC_VECTOR(7 DOWNTO 0)); 
END COMPONENT;

COMPONENT ULA is
    port(A, B: in STD_LOGIC_VECTOR(7 downto 0);
        S: in STD_LOGIC_VECTOR(2 downto 0);
        O: out STD_LOGIC_VECTOR(7 downto 0);
        C, Z: out STD_LOGIC);
END COMPONENT;

SIGNAL ULA_S, MUX_S, RP_DATA, RQ_DATA: STD_LOGIC_VECTOR(7 DOWNTO 0);


BEGIN 

MUX: MUX21_8 PORT MAP(R_DATA, ULA_S, MUX_SW, MUX_S);

BANCO: BANCO_REG168 PORT MAP(MUX_S, W_ADDR, RP_ADDR, RQ_ADDR, clr, CLK, W_WR, RP_RD, RQ_RD, RP_DATA, RQ_DATA);

ULAOP: ULA PORT MAP(RP_DATA, RQ_DATA, ULA_SW, ULA_S, ULA_CARRY, ULA_Z); 

S <= ULA_S;
W_DATA <= RP_DATA;

END CKT;