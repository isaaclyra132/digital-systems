library ieee;
use ieee.std_logic_1164.all;

ENTITY MUX16 IS
	PORT(EN, I0, I1, I2, I3, I4, I5, I6, I7, I8, I9, I10, I11, I12, I13, I14, I15: in STD_LOGIC;
		S: in STD_LOGIC_VECTOR(3 downto 0);
		O: out STD_LOGIC);
END MUX16;

ARCHITECTURE CKT OF MUX16 IS

BEGIN

	O <= EN AND ((I0 AND NOT S(3) AND NOT S(2) AND NOT S(1) AND NOT S(0)) 
	OR (I1 AND NOT S(3) AND NOT S(2) AND NOT S(1) AND S(0)) 
	OR (I2 AND NOT S(3) AND NOT S(2) AND S(1) AND NOT S(0))
	OR (I3 AND NOT S(3) AND NOT S(2) AND S(1) AND S(0)) 
	OR (I4 AND NOT S(3) AND S(2) AND NOT S(1) AND NOT S(0)) 
	OR (I5 AND NOT S(3) AND S(2) AND NOT S(1) AND S(0))
	OR (I6 AND NOT S(3) AND S(2) AND S(1) AND NOT S(0)) 
	OR (I7 AND NOT S(3) AND S(2) AND S(1) AND S(0)) 
	OR (I8 AND S(3) AND NOT S(2) AND NOT S(1) AND NOT S(0))
	OR (I9 AND S(3) AND NOT S(2) AND NOT S(1) AND S(0)) 
	OR (I10 AND S(3) AND NOT S(2) AND S(1) AND NOT S(0)) 
	OR (I11 AND S(3) AND NOT S(2) AND S(1) AND S(0))
	OR (I12 AND S(3) AND S(2) AND NOT S(1) AND NOT S(0))
	OR (I13 AND S(3) AND S(2) AND NOT S(1) AND S(0))
	OR (I14 AND S(3) AND S(2) AND S(1) AND NOT S(0))
	OR (I15 AND S(3) AND S(2) AND S(1) AND S(0)));

END CKT;